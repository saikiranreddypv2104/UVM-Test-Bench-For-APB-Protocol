`include "register_model.sv"
`include "bus_transaction.sv"
`include "transaction.sv"
`include "adapter.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "environment.sv"